module dynamic_op();
  int array[];
  initial begin
    array='{4,5,6,3,6,3};
    foreach(array[i])
      $display("array=%d",i,array[i]);
    $display("size of an array=%d",array.size());
    array.reverse();
    $display(array);
    array.sort();
    $display(array);
    array.rsort();
    $display(array);
    array.shuffle();
    $display(array);
    array.delete();
    $display("size of an array",array.size());
  end
endmodule
